** Profile: "SCHEMATIC1-sim2"  [ C:\USERS\LHLEE\APPDATA\ROAMING\SPB_DATA\CDSSETUP\WORKSPACE\PROJECTS\HW1\HW1-PSpiceFiles\SCHEMATIC1\sim2.sim ] 

** Creating circuit file "sim2.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\lhlee\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\24.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
